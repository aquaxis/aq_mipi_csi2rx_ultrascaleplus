module csi_rx_10b8b(
    input RST_M,
    input CLK,

    input [7:0]
);
endmodule
